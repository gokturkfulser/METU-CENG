`timescale 1ns / 1ps
module testbench_ic232;

	// write your code here
      
endmodule
