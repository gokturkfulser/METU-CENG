`timescale 1ns / 1ps
module testbench_numerator(
    );


endmodule
